`ifndef INCLUDE_TYPEDEF_COLLECTION_SV
`define INCLUDE_TYPEDEF_COLLECTION_SV

`define MEMSIZE 16
`define REGSIZE 8

typedef logic [`REGSIZE-1:0] DEFAULT_TYPE;

typedef enum logic [3:0] {
  RESET_STATE
  , FETCH_OPERATION
  , DECODE
  , FETCH_IMMEDIATE
  , FETCH_SRC
  , FETCH_SRC_IMM
  , FETCH_DST
  , FETCH_DST_IMM
  , EXECUTE
  , WRITE_REGISTER
  , WRITE_MEMORY
} STATE_TYPE;

typedef enum logic [3:0] {ADD, MOV, HLT, JMP} OPECODE_TYPE;

typedef enum logic [2:0] {REG_A, ADDRESS_REG_A, ADDRESS_IMM, IMM, UNUSED} OPERAND_TYPE;

typedef enum logic [3:0] {MEMORY_STAY, MEMORY_READ, MEMORY_WRITE} MEMORY_FLAG_TYPE;

`endif
